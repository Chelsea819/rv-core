/*************************************************************************
	> File Name: ysyx_23060025_counter.v
	> Author: Chelsea
	> Mail: 1938166340@qq.com 
	> Created Time: 2023年08月05日 星期六 22时12分23秒
 ************************************************************************/
// clock rstn waddr wdata wen wmask
`include "ysyx_23060025_define.v"
`include "ysyx_23060025_define_delay.v"
module ysyx_23060025_LSU #(parameter DATA_LEN = 32,ADDR_LEN = 32)(
	input								rstn			,
`ifdef DIFFTEST
	input								diff_skip_flag_i,
	output								diff_skip_flag_o,
`endif	
    input		                		wd_i		,
    input		                		clock			,
    input		[4:0]		            wreg_i		,
    input		[DATA_LEN - 1:0]		alu_result_i,
    input		                		mem_wen_i	,
	input		[DATA_LEN - 1:0]		mem_wdata_i	,
    input       [2:0]                   load_type_i , 
    input       [1:0]                   store_type_i, 
    input       [DATA_LEN - 1:0]        csr_wdata_i	,
    input       [11:0]       			csr_waddr_i	,
    input       [2:0]                   csr_type_i	,
	


	// exu_lsu
    input                                         exu_valid_i               ,
    output                                        lsu_ready_o               ,

    // lsu_wbu
    output                                        lsu_valid_o               ,
    input                                         wbu_ready_i               ,

	output                                        ebreak_flag_o               ,
    input                                         ebreak_flag_i               ,


    // input                               wb_ready_o  ,
    // output                              lsu_ready_o ,
    
    output	   	                		wd_o		,
    output	   	[4:0]		            wreg_o		,
	output     [DATA_LEN - 1:0]		    wdata_o,
    output      [DATA_LEN - 1:0]        csr_wdata_o	,
    output      [2:0]                   csr_type_o	,
	output       [11:0]        			csr_waddr_o	,
	// output                              memory_inst_o ,

    // AXI
    //Addr Read
	output		[ADDR_LEN - 1:0]		addr_r_addr_o,
	output		                		addr_r_valid_o,
	input		                		addr_r_ready_i,
	output		[2:0]                	addr_r_size_o,

	// Read data
	input		[DATA_LEN - 1:0]		r_data_i	,
	input		[1:0]					r_resp_i	,	// 读操作是否成功，存储器处理读写事物时可能会发生错误
	input		                		r_valid_i	,
	output		                		r_ready_o	,

	// Addr Write
	output		[ADDR_LEN - 1:0]		addr_w_addr_o,	// 写地址
	output		                		addr_w_valid_o,	// 主设备给出的地址和相关控制信号有效
	output		[2:0]                	addr_w_size_o,	// 主设备给出的地址和相关控制信号有效
	input		                		addr_w_ready_i, // 从设备已准备好接收地址和相关的控制信号

	// Write data
	output		[DATA_LEN - 1:0]		w_data_o	,	// 写出的数据
	output		[3:0]					w_strb_o	,	// wmask 	数据的字节选通，数据中每8bit对应这里的1bit
	output		                		w_valid_o	,	// 主设备给出的数据和字节选通信号有效
	input		                		w_ready_i	,	// 从设备已准备好接收数据选通信号

	// Backward
	input		[1:0]					bkwd_resp_i,	// 写回复信号，写操作是否成功
	input		                		bkwd_valid_i,	// 从设备给出的写回复信号是否有效
	output		                		bkwd_ready_o	// 主设备已准备好接收写回复信号
    
);	
    wire [31:0] mem_rdata;
	wire	 [DATA_LEN - 1:0]    mem_rdata_unaligned	;
	wire 		 				 aligned_store	;
    // reg  [7:0]  mem_rmask;
    wire        					mem_to_reg;
	wire	[3:0]					w_strb	;	// wmask 	数据的字节选通，数据中每8bit对应这里的1bit
	wire	[DATA_LEN - 1:0]		w_data	;	// wmask 	数据的字节选通，数据中每8bit对应这里的1bit

	assign ebreak_flag_o = ebreak_flag_i;
	assign csr_waddr_o = csr_waddr_i;
`ifdef DIFFTEST
	assign diff_skip_flag_o = diff_skip_flag_i;
`endif

	wire state_exe_valid = (con_state == STATE_WAIT_EXE_VALID);
	wire state_addr_pass = (con_state == LSU_WAIT_ADDR_PASS);
	wire state_data_load = (con_state == STATE_DATA_LOAD);
	reg			[1:0]			        	con_state	;
	reg			[1:0]			        	next_state	;
    parameter [1:0] STATE_WAIT_EXE_VALID = 2'b00, LSU_WAIT_ADDR_PASS = 2'b01, STATE_DATA_LOAD = 2'b11, LSU_WAIT_WB_READY = 2'b10;

    assign lsu_valid_o = (state_addr_pass && next_state == STATE_WAIT_EXE_VALID) 
						|| (state_data_load && next_state == STATE_WAIT_EXE_VALID) 
						|| next_state == LSU_WAIT_WB_READY;
    assign lsu_ready_o = state_exe_valid;

	// state trans
	always @(posedge clock ) begin
		if(rstn)
            con_state <= next_state;
		else 
			con_state <= STATE_WAIT_EXE_VALID;
	end


	// next_state
	always @(*) begin
		next_state = con_state;
		case(con_state) 
			STATE_WAIT_EXE_VALID: begin 
				if (exu_valid_i) begin
					next_state = LSU_WAIT_ADDR_PASS;
				end
			end
			LSU_WAIT_ADDR_PASS: begin 
				if(~(mem_to_reg | mem_wen_i)) begin 
					if(wbu_ready_i) begin
						next_state = STATE_WAIT_EXE_VALID;
					end else begin
						next_state = LSU_WAIT_WB_READY;
					end
                end else if (mem_to_reg & addr_r_ready_i) begin // read
					next_state = STATE_DATA_LOAD;
                end else if (mem_wen_i & addr_w_ready_i & w_ready_i & mem_wen_i) begin // read
					next_state = STATE_DATA_LOAD;
				end
			end
			STATE_DATA_LOAD: begin 
				if (r_valid_i | (~|bkwd_resp_i & bkwd_valid_i)) begin
					if(wbu_ready_i) begin
						next_state = STATE_WAIT_EXE_VALID;
					end else begin
						next_state = LSU_WAIT_WB_READY;
					end
					
				end
			end
            // 等待exu空闲，下LSU_WAIT_WB_READY个时钟周期传递信息
            LSU_WAIT_WB_READY: begin
				if (wbu_ready_i) begin
					next_state = STATE_WAIT_EXE_VALID;
				end
			end
            default: begin 
			end
		endcase
	end

	wire [31:0] r_data = r_data_i;


// delay test
`ifdef DELAY_TEST
	// random delay
	`ifdef RAN_DELAY
		reg				[3:0]		        	RANDOM_DELAY;
        reg				[3:0]		        	RANDOM_W_DATA_DELAY;
        wire			[3:0]		        	delay_num;
        wire			[3:0]		        	delay_num_w_data;

        ysyx_23060025_LFSR u_LFSR(
            .clock          ( clock          ),
            .rstn         ( rstn         ),
            .initial_var  ( 4'b1  		 ),
            .result       ( delay_num    )
        );
        ysyx_23060025_LFSR u_LFSR_w_data(
            .clock          ( clock          ),
            .rstn         ( rstn         ),
            .initial_var  ( 4'b1  		 ),
            .result       ( delay_num_w_data    )
        );
		
		always @(posedge clock ) begin
            if (~rstn) 
                RANDOM_DELAY <= 4'b1;
            else if((con_state == STATE_WAIT_EXE_VALID && next_state == LSU_WAIT_ADDR_PASS) || (con_state == LSU_WAIT_ADDR_PASS && next_state == LSU_WAIT_ADDR_PASS))
                RANDOM_DELAY <= delay_num;
        end

        always @(posedge clock ) begin
            if (~rstn) 
                RANDOM_W_DATA_DELAY <= 0;
            else if((con_state == STATE_WAIT_EXE_VALID && next_state == LSU_WAIT_ADDR_PASS))
                RANDOM_W_DATA_DELAY <= delay_num_w_data;
        end
	// fixed var delay
	`elsif VAR_DELAY
		// 当 RAN_DELAY 未定义，但 VAR_DELAY 被定义时，编译这段代码
        wire				[3:0]		        	RANDOM_DELAY;
        wire				[3:0]		        	RANDOM_W_DATA_DELAY;
		assign RANDOM_DELAY = `VAR_DELAY;
		assign RANDOM_W_DATA_DELAY = `VAR_W_DELAY;

	`endif

	reg			[3:0]		addr_r_valid_delay;
	reg			[3:0]		addr_w_valid_delay;
	reg			[3:0]		w_data_valid_delay;
	reg			[3:0]		r_ready_delay;
	reg			[3:0]		bkwd_ready_delay;

    assign addr_r_valid_o = (con_state == LSU_WAIT_ADDR_PASS) & mem_to_reg & rstn & (addr_r_valid_delay == RANDOM_DELAY); // addr valid and load inst
    assign r_ready_o = (con_state == LSU_WAIT_ADDR_PASS) & (r_ready_delay == RANDOM_DELAY);
    assign addr_w_valid_o = (con_state == LSU_WAIT_ADDR_PASS) & mem_wen_i & rstn & (addr_w_valid_delay == RANDOM_DELAY);  // addr valid and store inst
    assign w_valid_o = (con_state == LSU_WAIT_ADDR_PASS) & mem_wen_i & rstn & (w_data_valid_delay == RANDOM_W_DATA_DELAY);
    assign bkwd_ready_o = (con_state == LSU_WAIT_ADDR_PASS) & rstn & (bkwd_ready_delay == RANDOM_DELAY);

	// r addr delay
	always @(posedge clock ) begin
        if (next_state == LSU_WAIT_ADDR_PASS && (addr_r_valid_delay != RANDOM_DELAY || addr_r_valid_delay == 0))
			addr_r_valid_delay <= addr_r_valid_delay + 1;
		else if(next_state == LSU_WAIT_ADDR_PASS && addr_r_valid_delay == RANDOM_DELAY)
			addr_r_valid_delay <= addr_r_valid_delay;
		else 
			addr_r_valid_delay <= 4'b0;
	end
	always @(posedge clock ) begin
		if (next_state == LSU_WAIT_ADDR_PASS && (addr_w_valid_delay != RANDOM_DELAY || addr_w_valid_delay == 0))
			addr_w_valid_delay <= addr_w_valid_delay + 1;
        else if(next_state == LSU_WAIT_ADDR_PASS && addr_w_valid_delay == RANDOM_DELAY)
			addr_w_valid_delay <= addr_w_valid_delay;
		else  
			addr_w_valid_delay <= 4'b0;
	end
	always @(posedge clock ) begin
		if (next_state == LSU_WAIT_ADDR_PASS && (w_data_valid_delay != RANDOM_W_DATA_DELAY || w_data_valid_delay == 0))
			w_data_valid_delay <= w_data_valid_delay + 1;
        else if(next_state == LSU_WAIT_ADDR_PASS && w_data_valid_delay == RANDOM_W_DATA_DELAY)
			w_data_valid_delay <= w_data_valid_delay;
		else  
			w_data_valid_delay <= 4'b0;
	end

	always @(posedge clock ) begin
		if (next_state == LSU_WAIT_ADDR_PASS && (r_ready_delay != RANDOM_DELAY || r_ready_delay == 0)) 
			r_ready_delay <= r_ready_delay + 1;
		else if(next_state == LSU_WAIT_ADDR_PASS && r_ready_delay == RANDOM_DELAY)
			r_ready_delay <= r_ready_delay;
		else  
			r_ready_delay <= 4'b0;
	end
	always @(posedge clock ) begin
		if (next_state == LSU_WAIT_ADDR_PASS && (bkwd_ready_delay != RANDOM_DELAY || bkwd_ready_delay == 0)) 
			bkwd_ready_delay <= bkwd_ready_delay + 1;
		else if(next_state == LSU_WAIT_ADDR_PASS && bkwd_ready_delay == RANDOM_DELAY)
			bkwd_ready_delay <= bkwd_ready_delay;
		else 
			bkwd_ready_delay <= 4'b0;
	end
// no delay
`else
    assign addr_r_valid_o =  state_addr_pass & mem_to_reg; // addr valid and load inst
    assign r_ready_o = state_addr_pass | state_data_load;
    assign addr_w_valid_o = state_addr_pass & mem_wen_i;  // addr valid and store inst
    assign w_valid_o = state_addr_pass & mem_wen_i;
    assign bkwd_ready_o = state_addr_pass | state_data_load;

`endif

    // 写寄存器的信息
    wire		[DATA_LEN - 1:0]		    wdata       ;
    assign wdata = mem_to_reg ? mem_rdata : alu_result_i;

	assign addr_r_addr_o = alu_result_i;
	assign addr_w_addr_o = alu_result_i;
	assign w_strb = (store_type_i == `STORE_SB_8)? `AXI_W_STRB_8 :
                    (store_type_i == `STORE_SH_16) ? `AXI_W_STRB_16 :
                    (store_type_i == `STORE_SW_32) ? `AXI_W_STRB_32 : 
                    0;
	assign w_data = mem_wdata_i;
	
	assign addr_r_size_o = (load_type_i == `LOAD_LB_8)  ? `AXI_ADDR_SIZE_1 : 
							(load_type_i == `LOAD_LH_16) ? `AXI_ADDR_SIZE_2: 
							(load_type_i == `LOAD_LBU_8) ? `AXI_ADDR_SIZE_1: 
							(load_type_i == `LOAD_LHU_16) ? `AXI_ADDR_SIZE_2: 
							// (load_type_i == `LOAD_LW_32) ? `AXI_ADDR_SIZE_4: 
							`AXI_ADDR_SIZE_4;
							
	assign addr_w_size_o = (store_type_i == `STORE_SB_8)? `AXI_ADDR_SIZE_1 :
							(store_type_i == `STORE_SH_16) ? `AXI_ADDR_SIZE_2 :
							// (store_type_i == `STORE_SW_32) ? `AXI_ADDR_SIZE_4 : 
							`AXI_ADDR_SIZE_4;


`ifdef N_YOSYS_STA_CHECK
	// import "DPI-C" function void dtrace_func(int addr);
    // always @(*)
	// 	dtrace_func(addr_w_addr_o);
`ifdef PERFORMANCE_COUNTER
	import "DPI-C" function void lsu_p_counter_update();
	always @(posedge clock) begin
		if (state_exe_valid & next_state == LSU_WAIT_ADDR_PASS) begin
			lsu_p_counter_update();
		end
	end

	import "DPI-C" function void lsu_delay_counter_update();
	always @(posedge clock) begin
		if ((state_addr_pass & (mem_to_reg | mem_wen_i)) || state_data_load) begin
			lsu_delay_counter_update();
		end
	end
	`endif
`endif


	wire n_aligned_store = ~aligned_store;
	wire aligned = (alu_result_i[1:0] == 2'b00) | n_aligned_store;

	assign {w_strb_o, w_data_o} = aligned ? {w_strb, w_data} :
					alu_result_i[1:0] == 2'b01 ? {{w_strb[2:0], 1'b0}, {w_data[23:0], 8'b0}} :
					alu_result_i[1:0] == 2'b10 ? {{w_strb[1:0], 2'b0}, {w_data[15:0], 16'b0}} :
					alu_result_i[1:0] == 2'b11 ? {{w_strb[0], 3'b0}, {w_data[7:0], 24'b0}} : 0;

    assign wdata_o = wdata;


	// wire addr_unaligned = alu_result_i[1:0];

	wire addr_sram = (alu_result_i >= `DEVICE_SRAM_ADDR_L && alu_result_i <= `DEVICE_SRAM_ADDR_H);
	wire addr_flash = (alu_result_i >= `DEVICE_FLASH_ADDR_L && alu_result_i <= `DEVICE_FLASH_ADDR_H);
	wire addr_sdram = (alu_result_i >= `DEVICE_SDRAM_ADDR_L && alu_result_i <= `DEVICE_SDRAM_ADDR_H);
	wire addr_psram = (alu_result_i >= `DEVICE_PSRAM_ADDR_L && alu_result_i <= `DEVICE_PSRAM_ADDR_H);

	assign aligned_store = addr_sram | addr_flash | addr_sdram | addr_psram;

    assign  mem_to_reg = |load_type_i;

    // assign mem_ren_o = mem_to_reg;
    
    // load
	/*
		addr_unaligned--访存地址的后两位
		对于mem 地址0x80000010【0-3】-- 内容【00_01_02_03】
		PSRAM->CPU 00_01_02_03
		0x80000011 addr_unaligned[1:0] == 2'b01---- 【00_01_02_03】--[01_02_03_00]
		0x80000012 addr_unaligned[1:0] == 2'b10---- 【00_01_02_03】--[02_03_00_00]  
		0x80000013 addr_unaligned[1:0] == 2'b11---- 【00_01_02_03】--[03_00_00_00]
	*/

	assign mem_rdata_unaligned = (alu_result_i[1:0] == 2'b00 || n_aligned_store) ? {r_data} :
								alu_result_i[1:0] == 2'b01 ? {8'b0, {r_data[31:8]}} :
								alu_result_i[1:0] == 2'b10 ? {16'b0, {r_data[31:16]}} :
								alu_result_i[1:0] == 2'b11 ? {{24'b0, r_data[31:24]}} : 0;

								
    assign mem_rdata = (load_type_i == `LOAD_LB_8)  ? {{24{mem_rdata_unaligned[7]}}, mem_rdata_unaligned[7:0]} : 
                    (load_type_i == `LOAD_LH_16) ? {{16{mem_rdata_unaligned[15]}}, mem_rdata_unaligned[15:0]}: 
                    (load_type_i == `LOAD_LBU_8) ? {{24{1'b0}}, mem_rdata_unaligned[7:0]}: 
                    (load_type_i == `LOAD_LHU_16) ? {{16{1'b0}}, mem_rdata_unaligned[15:0]}: 
                    mem_rdata_unaligned;

    assign wd_o = wd_i;
    assign wreg_o = wreg_i;
    assign csr_wdata_o	     =     csr_wdata_i;  
    assign csr_type_o	     =     csr_type_i;  

endmodule

